module score_update (
  input wire [31:0] score,
  input wire hit_alien
);

//	always @* begin
//		if (hit_alien) begin
//			assign score = score + 5;
//		end
//	end
	
endmodule
